`define WAYS 3

extern void generate_test(int);



initial begin
    generate_test(`WAYS);    
end

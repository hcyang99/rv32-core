module dispatch(
    input ID_EX_PACKET [`WAYS-1: 0] id_packet_in;
    
    );